----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:29:33 12/01/2019 
-- Design Name: 
-- Module Name:    main_module - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity main_module is
	Port ( 
		var0 : in  STD_LOGIC;
		var1 : in  STD_LOGIC;
		var2 : in  STD_LOGIC;
		output0 : out STD_LOGIC;
		output1 : out STD_LOGIC;
		output2 : out STD_LOGIC
	);
end main_module;

architecture Behavioral of main_module is

begin


end Behavioral;

